//declaration of apb defines

`define ADDR_WIDTH 32

`define DATA_WIDTH 32

`define WAIT_READY 4
